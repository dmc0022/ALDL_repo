// hub75_phase1_pixel.v
// Phase 1: Single pixel moves across the panel, cycling R->G->B.
// Designed to drop into your existing top-level mux (same port list as hub75_uahlogo/hub75_gif).

module hub75_phase1_pixel #(
    parameter integer WIDTH          = 32,
    parameter integer ROWS_PER_GROUP = 16,   // 1/16 scan => 16 row addresses (top+bottom)
    parameter integer SHOW_TICKS     = 12000, // OE-on time per row (brightness / refresh tradeoff)
    parameter integer MOVE_FRAMES    = 20,    // move pixel every N full refreshes (speed)
    parameter         OE_ACTIVE_LOW  = 1      // most HUB75 panels: OE=0 enables output
)(
    input  wire       clk,
    input  wire       reset_n,

    output reg        r1,
    output reg        g1,
    output reg        b1,
    output reg        r2,
    output reg        g2,
    output reg        b2,

    output reg  [3:0] row_addr,
    output reg        clk_out,
    output reg        lat,
    output reg        oe
);

    // -------------------------
    // OE polarity helpers
    // -------------------------
    localparam OE_ON  = (OE_ACTIVE_LOW) ? 1'b0 : 1'b1;
    localparam OE_OFF = (OE_ACTIVE_LOW) ? 1'b1 : 1'b0;

    // -------------------------
    // Scan FSM: SHIFT -> LATCH -> SHOW
    // -------------------------
    localparam S_SHIFT = 2'd0;
    localparam S_LATCH = 2'd1;
    localparam S_SHOW  = 2'd2;

    reg [1:0] state;

    reg [5:0] col_idx;     // 0..31
    reg [3:0] row_idx;     // 0..15

    reg       shift_phase; // toggles to create a CLK pulse per column
    reg [15:0] show_cnt;   // enough bits for SHOW_TICKS

    // -------------------------
    // Moving pixel state (full 32x32)
    // -------------------------
    reg [5:0] pix_x;       // 0..31
    reg [5:0] pix_y;       // 0..31
    reg [1:0] color_sel;   // 0=R,1=G,2=B
    reg [15:0] move_frame_cnt;

    // Match logic for current scan row-pair

	 wire top_half = (pix_y < 6'd16);
	 wire bot_half = (pix_y >= 6'd16);
	 wire [3:0] pix_y_row = pix_y[3:0];

	 wire top_match = top_half && (row_idx == pix_y_row) && (col_idx == pix_x);
	 wire bot_match = bot_half && (row_idx == pix_y_row) && (col_idx == pix_x);

    // Color bits (1-bit channels for Phase 1 bring-up)
    wire c_r = (color_sel == 2'd0);
    wire c_g = (color_sel == 2'd1);
    wire c_b = (color_sel == 2'd2);

    // -------------------------
    // Sequential logic
    // -------------------------
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            // outputs
            r1 <= 0; g1 <= 0; b1 <= 0;
            r2 <= 0; g2 <= 0; b2 <= 0;
            row_addr <= 0;
            clk_out <= 0;
            lat <= 0;
            oe  <= OE_OFF;

            // fsm
            state <= S_SHIFT;
            col_idx <= 0;
            row_idx <= 0;
            shift_phase <= 0;
            show_cnt <= 0;

            // pixel motion
            pix_x <= 0;
            pix_y <= 0;
            color_sel <= 0;
            move_frame_cnt <= 0;

        end else begin
            // default “safe” values (overridden per-state)
            lat <= 1'b0;

            // Keep row_addr updated to current scan row
            row_addr <= row_idx;

            case (state)

                // ---------------------------------
                // SHIFT: present RGB data + pulse CLK for each column
                // ---------------------------------
                S_SHIFT: begin
                    oe <= OE_OFF;     // blank while shifting
                    clk_out <= 1'b0;  // default low

                    // Only drive pixel data on the setup half-cycle
                    if (shift_phase == 1'b0) begin
                        // Drive RGB for this column and current row-pair
                        r1 <= top_match ? c_r : 1'b0;
                        g1 <= top_match ? c_g : 1'b0;
                        b1 <= top_match ? c_b : 1'b0;

                        r2 <= bot_match ? c_r : 1'b0;
                        g2 <= bot_match ? c_g : 1'b0;
                        b2 <= bot_match ? c_b : 1'b0;

                        // Next cycle will be the rising edge pulse
                        shift_phase <= 1'b1;

                    end else begin
                        // Pulse panel CLK (rising edge shifts current column)
                        clk_out <= 1'b1;

                        // Finish this column; advance column counter
                        shift_phase <= 1'b0;

                        if (col_idx == WIDTH-1) begin
                            col_idx <= 0;
                            state   <= S_LATCH;
                        end else begin
                            col_idx <= col_idx + 1'b1;
                        end
                    end
                end

                // ---------------------------------
                // LATCH: commit shifted row data
                // ---------------------------------
                S_LATCH: begin
                    oe      <= OE_OFF; // still blank
                    clk_out <= 1'b0;
                    lat     <= 1'b1;   // 1-cycle latch pulse
                    show_cnt <= 0;
                    state   <= S_SHOW;
                end

                // ---------------------------------
                // SHOW: enable LEDs for SHOW_TICKS
                // ---------------------------------
                S_SHOW: begin
                    clk_out <= 1'b0;
                    oe      <= OE_ON;

                    if (show_cnt == SHOW_TICKS-1) begin
                        oe <= OE_OFF;      // blank before next row shift
                        show_cnt <= 0;

                        // Advance row
                        if (row_idx == ROWS_PER_GROUP-1) begin
                            row_idx <= 0;

                            // End of full refresh frame -> update move timer
                            if (move_frame_cnt == MOVE_FRAMES-1) begin
                                move_frame_cnt <= 0;

                                // Move pixel across full 32x32 (row-major)
                                if (pix_x == WIDTH-1) begin
                                    pix_x <= 0;
                                    if (pix_y == (2*ROWS_PER_GROUP)-1)
                                        pix_y <= 0;
                                    else
                                        pix_y <= pix_y + 1'b1;
                                end else begin
                                    pix_x <= pix_x + 1'b1;
                                end

                                // Cycle color R -> G -> B -> R ...
                                if (color_sel == 2'd2)
                                    color_sel <= 2'd0;
                                else
                                    color_sel <= color_sel + 1'b1;

                            end else begin
                                move_frame_cnt <= move_frame_cnt + 1'b1;
                            end

                        end else begin
                            row_idx <= row_idx + 1'b1;
                        end

                        // Back to shifting next row
                        state <= S_SHIFT;

                    end else begin
                        show_cnt <= show_cnt + 1'b1;
                    end
                end

                default: begin
                    state <= S_SHIFT;
                end
            endcase
        end
    end

endmodule
